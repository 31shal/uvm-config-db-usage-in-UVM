interface mem_if(input clk, input reset);
logic [7:0]addr;
logic rden;
logic wren;
logic [31:0]read_data;
logic [31:0]write_data;
logic valid;  
endinterface: mem_if
